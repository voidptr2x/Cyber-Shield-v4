module utils

pub fn place_text(position []string, text string)
{
	print("")
}