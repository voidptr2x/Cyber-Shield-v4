module tools

pub struct System
{
	pub mut:
		con			Connection
		os			OS
		hdw			Hardware
		ui_mode		bool
}